* E:\Dropbox\JERRYL WORK\LT Spice Files\N-channel_MOSFET_L=5,W=10\N-channel_MOSFET.cir
.end
